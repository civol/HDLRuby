/* Description of an 8-bit data 8-bit address rom. */

module rom(en,rwb,addr,data);

    input[7:0]       addr;
    output reg [7:0] data;

    reg [7:0] content[0:255];

    always @ (*)
    begin
        case(addr)
            0: data <= 0;
            1: data <= 1;
            2: data <= 2;
            3: data <= 3;
            4: data <= 4;
            5: data <= 5;
            6: data <= 6;
            7: data <= 7;
            8: data <= 8;
            9: data <= 9;
            10: data <= 10;
            11: data <= 11;
            12: data <= 12;
            13: data <= 13;
            14: data <= 14;
            15: data <= 15;
            16: data <= 16;
            17: data <= 17;
            18: data <= 18;
            19: data <= 19;
            20: data <= 20;
            21: data <= 21;
            22: data <= 22;
            23: data <= 23;
            24: data <= 16;
            25: data <= 25;
            26: data <= 26;
            27: data <= 27;
            28: data <= 28;
            29: data <= 29;
            30: data <= 30;
            31: data <= 31;
            32: data <= 32;
            33: data <= 33;
            34: data <= 34;
            35: data <= 35;
            36: data <= 36;
            37: data <= 37;
            38: data <= 38;
            39: data <= 39;
            40: data <= 40;
            41: data <= 41;
            42: data <= 42;
            43: data <= 43;
            44: data <= 44;
            45: data <= 45;
            46: data <= 46;
            47: data <= 47;
            48: data <= 48;
            49: data <= 49;
            50: data <= 50;
            51: data <= 51;
            52: data <= 52;
            53: data <= 53;
            54: data <= 54;
            55: data <= 55;
            56: data <= 48;
            57: data <= 57;
            58: data <= 58;
            59: data <= 59;
            60: data <= 60;
            61: data <= 61;
            62: data <= 62;
            63: data <= 63;
            64: data <= 64;
            65: data <= 65;
            66: data <= 66;
            67: data <= 67;
            68: data <= 68;
            69: data <= 69;
            70: data <= 70;
            71: data <= 71;
            72: data <= 72;
            73: data <= 73;
            74: data <= 74;
            75: data <= 75;
            76: data <= 76;
            77: data <= 77;
            78: data <= 78;
            79: data <= 79;
            80: data <= 80;
            81: data <= 81;
            82: data <= 82;
            83: data <= 83;
            84: data <= 84;
            85: data <= 85;
            86: data <= 86;
            87: data <= 87;
            88: data <= 80;
            89: data <= 89;
            90: data <= 90;
            91: data <= 91;
            92: data <= 92;
            93: data <= 93;
            94: data <= 94;
            95: data <= 95;
            96: data <= 96;
            97: data <= 97;
            98: data <= 98;
            99: data <= 99;
            100: data <= 100;
            101: data <= 101;
            102: data <= 102;
            103: data <= 103;
            104: data <= 104;
            105: data <= 105;
            106: data <= 106;
            107: data <= 107;
            108: data <= 108;
            109: data <= 109;
            110: data <= 110;
            111: data <= 111;
            112: data <= 112;
            113: data <= 113;
            114: data <= 114;
            115: data <= 115;
            116: data <= 116;
            117: data <= 117;
            118: data <= 118;
            119: data <= 119;
            120: data <= 112;
            121: data <= 121;
            122: data <= 122;
            123: data <= 123;
            124: data <= 124;
            125: data <= 125;
            126: data <= 126;
            127: data <= 127;
            128: data <= 128;
            129: data <= 129;
            130: data <= 130;
            131: data <= 131;
            132: data <= 132;
            133: data <= 133;
            134: data <= 134;
            135: data <= 135;
            136: data <= 136;
            137: data <= 137;
            138: data <= 138;
            139: data <= 139;
            140: data <= 140;
            141: data <= 141;
            142: data <= 142;
            143: data <= 143;
            144: data <= 144;
            145: data <= 145;
            146: data <= 146;
            147: data <= 147;
            148: data <= 148;
            149: data <= 149;
            150: data <= 150;
            151: data <= 151;
            152: data <= 144;
            153: data <= 153;
            154: data <= 154;
            155: data <= 155;
            156: data <= 156;
            157: data <= 157;
            158: data <= 158;
            159: data <= 159;
            160: data <= 160;
            161: data <= 161;
            162: data <= 162;
            163: data <= 163;
            164: data <= 164;
            165: data <= 165;
            166: data <= 166;
            167: data <= 167;
            168: data <= 168;
            169: data <= 169;
            170: data <= 170;
            171: data <= 171;
            172: data <= 172;
            173: data <= 173;
            174: data <= 174;
            175: data <= 175;
            176: data <= 176;
            177: data <= 177;
            178: data <= 178;
            179: data <= 179;
            180: data <= 180;
            181: data <= 181;
            182: data <= 182;
            183: data <= 183;
            184: data <= 176;
            185: data <= 185;
            186: data <= 186;
            187: data <= 187;
            188: data <= 188;
            189: data <= 189;
            190: data <= 190;
            191: data <= 191;
            192: data <= 192;
            193: data <= 193;
            194: data <= 194;
            195: data <= 195;
            196: data <= 196;
            197: data <= 197;
            198: data <= 198;
            199: data <= 199;
            200: data <= 200;
            201: data <= 201;
            202: data <= 202;
            203: data <= 203;
            204: data <= 204;
            205: data <= 205;
            206: data <= 206;
            207: data <= 207;
            208: data <= 208;
            209: data <= 209;
            210: data <= 210;
            211: data <= 211;
            212: data <= 212;
            213: data <= 213;
            214: data <= 214;
            215: data <= 215;
            216: data <= 208;
            217: data <= 217;
            218: data <= 218;
            219: data <= 219;
            220: data <= 220;
            221: data <= 221;
            222: data <= 222;
            223: data <= 223;
            224: data <= 224;
            225: data <= 225;
            226: data <= 226;
            227: data <= 227;
            228: data <= 228;
            229: data <= 229;
            230: data <= 230;
            231: data <= 231;
            232: data <= 232;
            233: data <= 233;
            234: data <= 234;
            235: data <= 235;
            236: data <= 236;
            237: data <= 237;
            238: data <= 238;
            239: data <= 239;
            240: data <= 240;
            241: data <= 241;
            242: data <= 242;
            243: data <= 243;
            244: data <= 244;
            245: data <= 245;
            246: data <= 246;
            247: data <= 247;
            248: data <= 240;
            249: data <= 249;
            250: data <= 250;
            251: data <= 251;
            252: data <= 252;
            253: data <= 253;
            254: data <= 254;
            255: data <= 255;
        endcase
    end

endmodule
